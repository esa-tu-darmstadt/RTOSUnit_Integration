module cv32e40p_tb_top (
    // Clock and Reset
    input logic clk_i,
    input logic rst_ni,

    input logic pulp_clock_en_i,  // PULP clock enable (only used if COREV_CLUSTER = 1)
    input logic scan_cg_en_i,  // Enable all clock gates for testing

    // Core ID, Cluster ID, debug mode halt address and boot address are considered more or less static
    input logic [31:0] boot_addr_i,
    input logic [31:0] mtvec_addr_i,
    input logic [31:0] dm_halt_addr_i,
    input logic [31:0] hart_id_i,
    input logic [31:0] dm_exception_addr_i,

    // Instruction memory interface
    output logic        instr_req_o,
    input  logic        instr_gnt_i,
    input  logic        instr_rvalid_i,
    output logic [31:0] instr_addr_o,
    input  logic [31:0] instr_rdata_i,

    // Data memory interface
    output logic        data_req_o,
    input  logic        data_gnt_i,
    input  logic        data_rvalid_i,
    output logic        data_we_o,
    output logic [ 3:0] data_be_o,
    output logic [31:0] data_addr_o,
    output logic [31:0] data_wdata_o,
    input  logic [31:0] data_rdata_i,

    // Interrupt inputs
    input  logic [31:0] irq_i,  // CLINT interrupts + CLINT extension interrupts
    output logic        irq_ack_o,
    output logic [ 4:0] irq_id_o,

    // Debug Interface
    input  logic debug_req_i,
    output logic debug_havereset_o,
    output logic debug_running_o,
    output logic debug_halted_o,

    // CPU Control Signals
    input  logic fetch_enable_i,
    output logic core_sleep_o
);

// latch response from OBI
logic        data_rvalid_d;
logic [31:0] data_rdata_d;

always_ff @(posedge clk_i) begin
    data_rvalid_d <= data_rvalid_i;
    data_rdata_d <= data_rdata_i;
end

// Register Read Logic
logic [4:0] reg_read_addr_cold_u_to_c;          // reg_read_addr_cold
logic [31:0] reg_read_data_cold_data_c_to_u;    // reg_read_data_cold_data

// Register Write Logic
logic [36:0] reg_write_cold_u_to_c;             // reg_write_cold
logic RDY_reg_write_cold_u_to_c;                // RDY_reg_write_cold

// Cold Registers Logic
logic [927:0] cold_regs_in_c_to_u;              // cold_regs_in

// Hot Register Write Logic
logic [11:0] reg_hot_write_trace_addrs_c_to_u;    // reg_hot_write_trace_addr

// Mstatus and Mepc Logic
logic [31:0] mstatus_out_u_to_c;                // mstatus_out
logic [31:0] mepc_out_u_to_c;                   // mepc_out

// Bank Switching Logic
logic switch_bank_o_u_to_c;                     // switch_bank_o

// Mret Logic
logic EN_mret_c_to_u;                           // EN_mret
logic mret_u_to_c;                              // mret
logic RDY_mret_u_to_c;                          // RDY_mret

// CSR Write Logic
logic write_csrs_u_to_c;                        // write_csrs

// Trap Logic
logic [31:0] trap_mstatus_c_to_u;               // trap_mstatus
logic [31:0] trap_mepc_c_to_u;                  // trap_mepc
logic [31:0] trap_mcause_c_to_u;                // trap_mcause
logic EN_trap_c_to_u;                           // EN_trap
logic RDY_trap_u_to_c;                          // RDY_trap

// Custom Instruction Logic
logic [2:0] custom_inst_funct3_c_to_u;          // custom_inst_funct3
logic [31:0] custom_inst_id_c_to_u;             // custom_inst_id
logic [31:0] custom_inst_prio_c_to_u;           // custom_inst_prio
logic EN_custom_inst_c_to_u;                    // EN_custom_inst
logic [32:0] custom_inst_u_to_c;                // custom_inst
logic RDY_custom_inst_u_to_c;                   // RDY_custom_inst

// memory bus arbitration
logic        data_req_c;
logic        data_gnt_c;
logic        data_rvalid_c;
logic        data_we_c;
logic [ 3:0] data_be_c;
logic [31:0] data_addr_c;
logic [31:0] data_wdata_c;
logic [31:0] data_rdata_c;

assign data_gnt_c = data_gnt_i;

logic [64:0] ctx_mem_access;
logic        EN_ctx_mem_access;
logic        RDY_ctx_mem_access;

// internal signals for RTOSUnit memory iface
logic        ctx_mem_wr_en;
logic [31:0] ctx_mem_addr;
logic [31:0] ctx_mem_wr_data;
logic ctx_mem_rd_rq_valid;

// request source tracking
logic [1:0] rq_ptr;
logic [1:0] rs_ptr;
logic [2:0] src_arr [3:0];

logic ctx_mem_rd_resp_valid;
logic [31:0] ctx_mem_rd_data;

// store source of a request
always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
        rq_ptr <= 0;
        rs_ptr <= 0;
    end else begin
        src_arr[rq_ptr] <= {data_req_c, ctx_mem_wr_en && EN_ctx_mem_access, EN_ctx_mem_access && ~ctx_mem_wr_en};
        if (data_req_c | EN_ctx_mem_access) begin
            rq_ptr <= rq_ptr + 1;
        end
    end
end

// distribute incoming reads
always_comb begin
    data_rdata_c = data_rdata_d;
    ctx_mem_rd_data = data_rdata_d;

    data_rvalid_c         = data_rvalid_d & src_arr[rs_ptr][2];
    ctx_mem_rd_resp_valid = data_rvalid_d & src_arr[rs_ptr][0];
end

// advance response destination pointer
always_ff @(posedge clk_i) begin
    if (rst_ni && data_rvalid_d) rs_ptr <= rs_ptr + 1;
end

// arbitrate memory bus between CPU and RTOSUNIT
assign EN_ctx_mem_access = ~data_req_c & RDY_ctx_mem_access;
assign ctx_mem_addr      = ctx_mem_access[64:33];
assign ctx_mem_wr_data   = ctx_mem_access[32:1];
assign ctx_mem_wr_en     = ctx_mem_access[0];

// build output signals for memory bus
always_comb begin
    data_req_o   = data_req_c | EN_ctx_mem_access;

    data_we_o    = data_req_c ?    data_we_c  :  ctx_mem_wr_en;
    data_be_o    = data_req_c ?    data_be_c  :  'hf;
    data_addr_o  = data_req_c ?  data_addr_c  :  ctx_mem_addr;
    data_wdata_o = data_req_c ? data_wdata_c  :  ctx_mem_wr_data;
end

// write request separation
logic [4:0] reg_write_cold_addr;
logic [31:0] reg_write_cold_data;
assign reg_write_cold_addr = reg_write_cold_u_to_c[36:32];
assign reg_write_cold_data = reg_write_cold_u_to_c[31:0];

cv32e40p_core #(
    .FPU                      ( 0 ),
    .FPU_ADDMUL_LAT           ( 0 ),
    .FPU_OTHERS_LAT           ( 0 ),
    .ZFINX                    ( 0 ),
    .COREV_PULP               ( 0 ),
    .COREV_CLUSTER            ( 0 ),
    .NUM_MHPMCOUNTERS         ( 1 )
) u_core (
    // Clock and reset
    .rst_ni                   (rst_ni),
    .clk_i                    (clk_i),
    .scan_cg_en_i             (scan_cg_en_i),

    // Special control signals
    .fetch_enable_i           (fetch_enable_i),
    .pulp_clock_en_i          (pulp_clock_en_i),
    .core_sleep_o             (core_sleep_o),

    // Configuration
    .boot_addr_i              (boot_addr_i),
    .mtvec_addr_i             (mtvec_addr_i),
    .dm_halt_addr_i           (dm_halt_addr_i),
    .dm_exception_addr_i      (dm_exception_addr_i),
    .hart_id_i                (hart_id_i),

    // Instruction memory interface
    .instr_addr_o             (instr_addr_o),
    .instr_req_o              (instr_req_o),
    .instr_gnt_i              (instr_gnt_i),
    .instr_rvalid_i           (instr_rvalid_i),
    .instr_rdata_i            (instr_rdata_i),

    // Data memory interface
    .data_addr_o              (data_addr_c),
    .data_req_o               (data_req_c),
    .data_gnt_i               (data_gnt_c),
    .data_we_o                (data_we_c),
    .data_be_o                (data_be_c),
    .data_wdata_o             (data_wdata_c),
    .data_rvalid_i            (data_rvalid_c),
    .data_rdata_i             (data_rdata_c),

     // Interrupt interface
    .irq_i                    (irq_i),
    .irq_ack_o                (irq_ack_o),
    .irq_id_o                 (irq_id_o),

    // Debug interface
    .debug_req_i              (debug_req_i),
    .debug_havereset_o        (debug_havereset_o),
    .debug_running_o          (debug_running_o),
    .debug_halted_o           (debug_halted_o),

    // ctx operations
    .ctx_en_op_o(EN_custom_inst_c_to_u),
    .ctx_op_funct3_o(custom_inst_funct3_c_to_u),
    .ctx_rs1_id_o(custom_inst_id_c_to_u),
    .ctx_rs2_prio_o(custom_inst_prio_c_to_u),
    .ctx_rd_write_data_i(custom_inst_u_to_c),
    .ctx_mret_o(EN_mret_c_to_u),
    .ctx_trap_o(EN_trap_c_to_u),

    // ctx reg access
    .reg_read_addr_cold_i(reg_read_addr_cold_u_to_c),
    .reg_read_data_cold_data_o(reg_read_data_cold_data_c_to_u),

    .reg_write_addr_cold_i(reg_write_cold_addr),
    .reg_write_data_cold_data_i(reg_write_cold_data),
    .reg_write_we_cold_i(RDY_reg_write_cold_u_to_c),

    // ctx stuff
    .ctx_mcause_o(trap_mcause_c_to_u),
    .ctx_mstatus_o(trap_mstatus_c_to_u),
    .ctx_mepc_o(trap_mepc_c_to_u),
    .ctx_switch_bank_i(switch_bank_o_u_to_c),

    .ctx_csr_wr_we_i(write_csrs_u_to_c),
    .ctx_csr_wr_mepc_i(mepc_out_u_to_c),
    .ctx_csr_wr_mstatus_i(mstatus_out_u_to_c),

    .ctx_stall_mret_i(~RDY_mret_u_to_c),

    .ctx_reg_hot_write_trace_o(reg_hot_write_trace_addrs_c_to_u),

    .apu_busy_o    (),
    .apu_req_o     (),
    .apu_gnt_i     (0),
    .apu_operands_o(),
    .apu_op_o      (),
    .apu_flags_o   (),
    .apu_rvalid_i  (0),
    .apu_result_i  (0),
    .apu_flags_i   (0)
);

// Instantiate mkRTOSUnitSynth
mkRTOSUnitSynth u_mkRTOSUnitSynth (
    .CLK                        (clk_i),                      // Clock input
    .RST_N                      (rst_ni),                    // Reset input

    // Register Read Logic
    .reg_read_addr_cold         (reg_read_addr_cold_u_to_c), // reg_read_addr_cold
    .reg_read_data_cold_data    (reg_read_data_cold_data_c_to_u), // reg_read_data_cold_data

    // Register Write Logic
    .EN_reg_write_cold          (RDY_reg_write_cold_u_to_c), // EN_reg_write_cold
    .reg_write_cold             (reg_write_cold_u_to_c),    // reg_write_cold
    .RDY_reg_write_cold         (RDY_reg_write_cold_u_to_c), // RDY_reg_write_cold

    // Cold Registers Logic
    .cold_regs_in               (cold_regs_in_c_to_u),      // cold_regs_in

    // Hot Register Write Logic
    .reg_hot_write_trace_addrs   (reg_hot_write_trace_addrs_c_to_u), // reg_hot_write_trace_addr

    // Memory Write Logic
    /*.EN_mem_wr                  (EN_mem_wr_c_to_u),         // EN_mem_wr
    .mem_wr                     (mem_wr_u_to_c),            // mem_wr
    .RDY_mem_wr                 (RDY_mem_wr_u_to_c),        // RDY_mem_wr*/

    /*// Memory Read Address Logic
    .EN_mem_rd_addr             (ctx_mem_rd_rq_valid),    // EN_mem_rd_addr
    .mem_rd_addr                (ctx_mem_rd_rq_addr),       // mem_rd_addr
    .RDY_mem_rd_addr            (RDY_mem_rd_addr_u_to_c),   // RDY_mem_rd_addr*/

    // Memory Read Data Logic
    .mem_rd_data_d              (ctx_mem_rd_data),     // mem_rd_data_d
    .EN_mem_rd_data             (ctx_mem_rd_resp_valid),    // EN_mem_rd_data

    .mem_access                 (ctx_mem_access),
    .EN_mem_access              (EN_ctx_mem_access),
    .RDY_mem_access             (RDY_ctx_mem_access),

    // Mstatus and Mepc Logic
    .mstatus_out                (mstatus_out_u_to_c),       // mstatus_out
    .mepc_out                   (mepc_out_u_to_c),          // mepc_out

    // Bank Switching Logic
    .switch_bank_o              (switch_bank_o_u_to_c),     // switch_bank_o

    // Mret Logic
    .EN_mret                    (EN_mret_c_to_u),           // EN_mret
    .mret                       (mret_u_to_c),              // mret
    .RDY_mret                   (RDY_mret_u_to_c),          // RDY_mret

    // CSR Write Logic
    .write_csrs                 (write_csrs_u_to_c),        // write_csrs

    // Trap Logic
    .trap_mstatus               (trap_mstatus_c_to_u),      // trap_mstatus
    .trap_mepc                  (trap_mepc_c_to_u),         // trap_mepc
    .trap_mcause                (trap_mcause_c_to_u),       // trap_mcause
    .EN_trap                    (EN_trap_c_to_u),           // EN_trap
    .RDY_trap                   (RDY_trap_u_to_c),          // RDY_trap

    // Custom Instruction Logic
    .custom_inst_funct3         (custom_inst_funct3_c_to_u),// custom_inst_funct3
    .custom_inst_id             (custom_inst_id_c_to_u),    // custom_inst_id
    .custom_inst_prio           (custom_inst_prio_c_to_u),  // custom_inst_prio
    .EN_custom_inst             (EN_custom_inst_c_to_u),    // EN_custom_inst
    .custom_inst                (custom_inst_u_to_c),       // custom_inst
    .RDY_custom_inst            (RDY_custom_inst_u_to_c)    // RDY_custom_inst
);



endmodule
