// Copyright 2017-2019 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Author: Florian Zaruba, ETH Zurich
// Date: 19.03.2017
// Description: CVA6 Top-level module

`include "rvfi_types.svh"
`include "cvxif_types.svh"

module cva6_ariane_wrapper import ariane_pkg::*; #(
    // CVA6 config
    parameter config_pkg::cva6_cfg_t CVA6Cfg = build_config_pkg::build_config(
        cva6_config_pkg::cva6_cfg
    ),

    // RVFI PROBES
    parameter type rvfi_probes_instr_t = `RVFI_PROBES_INSTR_T(CVA6Cfg),
    parameter type rvfi_probes_csr_t = `RVFI_PROBES_CSR_T(CVA6Cfg),
    parameter type rvfi_probes_t = struct packed {
      logic csr;
      rvfi_probes_instr_t instr;
    },

    // branchpredict scoreboard entry
    // this is the struct which we will inject into the pipeline to guide the various
    // units towards the correct branch decision and resolve
    localparam type branchpredict_sbe_t = struct packed {
      cf_t                     cf;               // type of control flow prediction
      logic [CVA6Cfg.VLEN-1:0] predict_address;  // target address at which to jump, or not
    },

    localparam type exception_t = struct packed {
      logic [CVA6Cfg.XLEN-1:0] cause;  // cause of exception
      logic [CVA6Cfg.XLEN-1:0] tval;  // additional information of causing exception (e.g.: instruction causing it),
      // address of LD/ST fault
      logic [CVA6Cfg.GPLEN-1:0] tval2;  // additional information when the causing exception in a guest exception
      logic [31:0] tinst;  // transformed instruction information
      logic gva;  // signals when a guest virtual address is written to tval
      logic valid;
    },

    // cache request ports
    // I$ address translation requests
    localparam type icache_areq_t = struct packed {
      logic                    fetch_valid;      // address translation valid
      logic [CVA6Cfg.PLEN-1:0] fetch_paddr;      // physical address in
      exception_t              fetch_exception;  // exception occurred during fetch
    },
    localparam type icache_arsp_t = struct packed {
      logic                    fetch_req;    // address translation request
      logic [CVA6Cfg.VLEN-1:0] fetch_vaddr;  // virtual address out
    },

    // I$ data requests
    localparam type icache_dreq_t = struct packed {
      logic                    req;      // we request a new word
      logic                    kill_s1;  // kill the current request
      logic                    kill_s2;  // kill the last request
      logic                    spec;     // request is speculative
      logic [CVA6Cfg.VLEN-1:0] vaddr;    // 1st cycle: 12 bit index is taken for lookup
    },
    localparam type icache_drsp_t = struct packed {
      logic                                ready;  // icache is ready
      logic                                valid;  // signals a valid read
      logic [CVA6Cfg.FETCH_WIDTH-1:0]      data;   // 2+ cycle out: tag
      logic [CVA6Cfg.FETCH_USER_WIDTH-1:0] user;   // User bits
      logic [CVA6Cfg.VLEN-1:0]             vaddr;  // virtual address out
      exception_t                          ex;     // we've encountered an exception
    },

    // IF/ID Stage
    // store the decompressed instruction
    localparam type fetch_entry_t = struct packed {
      logic [CVA6Cfg.VLEN-1:0] address;  // the address of the instructions from below
      logic [31:0] instruction;  // instruction word
      branchpredict_sbe_t     branch_predict; // this field contains branch prediction information regarding the forward branch path
      exception_t             ex;             // this field contains exceptions which might have happened earlier, e.g.: fetch exceptions
    },

    // ID/EX/WB Stage
    localparam type scoreboard_entry_t = struct packed {
      logic [CVA6Cfg.VLEN-1:0] pc;  // PC of instruction
      logic [CVA6Cfg.TRANS_ID_BITS-1:0] trans_id;      // this can potentially be simplified, we could index the scoreboard entry
      // with the transaction id in any case make the width more generic
      fu_t fu;  // functional unit to use
      fu_op op;  // operation to perform in each functional unit
      logic [REG_ADDR_SIZE-1:0] rs1;  // register source address 1
      logic [REG_ADDR_SIZE-1:0] rs2;  // register source address 2
      logic [REG_ADDR_SIZE-1:0] rd;  // register destination address
      logic [CVA6Cfg.XLEN-1:0] result;  // for unfinished instructions this field also holds the immediate,
      // for unfinished floating-point that are partly encoded in rs2, this field also holds rs2
      // for unfinished floating-point fused operations (FMADD, FMSUB, FNMADD, FNMSUB)
      // this field holds the address of the third operand from the floating-point register file
      logic valid;  // is the result valid
      logic use_imm;  // should we use the immediate as operand b?
      logic use_zimm;  // use zimm as operand a
      logic use_pc;  // set if we need to use the PC as operand a, PC from exception
      exception_t ex;  // exception has occurred
      branchpredict_sbe_t bp;  // branch predict scoreboard data structure
      logic                     is_compressed; // signals a compressed instructions, we need this information at the commit stage if
                                               // we want jump accordingly e.g.: +4, +2
      logic is_macro_instr;  // is an instruction executed as predefined sequence of instructions called macro definition
      logic is_last_macro_instr;  // is last decoded 32bit instruction of macro definition
      logic is_double_rd_macro_instr;  // is double move decoded 32bit instruction of macro definition
      logic vfp;  // is this a vector floating-point instruction?
    },

    // branch-predict
    // this is the struct we get back from ex stage and we will use it to update
    // all the necessary data structures
    // bp_resolve_t
    localparam type bp_resolve_t = struct packed {
      logic                    valid;           // prediction with all its values is valid
      logic [CVA6Cfg.VLEN-1:0] pc;              // PC of predict or mis-predict
      logic [CVA6Cfg.VLEN-1:0] target_address;  // target address at which to jump, or not
      logic                    is_mispredict;   // set if this was a mis-predict
      logic                    is_taken;        // branch is taken
      cf_t                     cf_type;         // Type of control flow change
    },

    // All information needed to determine whether we need to associate an interrupt
    // with the corresponding instruction or not.
    localparam type irq_ctrl_t = struct packed {
      logic [CVA6Cfg.XLEN-1:0] mie;
      logic [CVA6Cfg.XLEN-1:0] mip;
      logic [CVA6Cfg.XLEN-1:0] mideleg;
      logic [CVA6Cfg.XLEN-1:0] hideleg;
      logic                    sie;
      logic                    global_enable;
    },

    localparam type lsu_ctrl_t = struct packed {
      `ifdef SCAIEV_MEM
      logic 							rdMem_ISAX;
      `endif
      logic                             valid;
      logic [CVA6Cfg.VLEN-1:0]          vaddr;
      logic [31:0]                      tinst;
      logic                             hs_ld_st_inst;
      logic                             hlvx_inst;
      logic                             overflow;
      logic                             g_overflow;
      logic [CVA6Cfg.XLEN-1:0]          data;
      logic [(CVA6Cfg.XLEN/8)-1:0]      be;
      fu_t                              fu;
      fu_op                             operation;
      logic [CVA6Cfg.TRANS_ID_BITS-1:0] trans_id;
    },

    localparam type fu_data_t = struct packed {
      fu_t                              fu;
      fu_op                             operation;
      logic [CVA6Cfg.XLEN-1:0]          operand_a;
      logic [CVA6Cfg.XLEN-1:0]          operand_b;
      logic [CVA6Cfg.XLEN-1:0]          imm;
      logic [CVA6Cfg.TRANS_ID_BITS-1:0] trans_id;
    },

    localparam type icache_req_t = struct packed {
      logic [CVA6Cfg.ICACHE_SET_ASSOC_WIDTH-1:0] way;  // way to replace
      logic [CVA6Cfg.PLEN-1:0] paddr;  // physical address
      logic nc;  // noncacheable
      logic [CVA6Cfg.MEM_TID_WIDTH-1:0] tid;  // threadi id (used as transaction id in Ariane)
    },
    localparam type icache_rtrn_t = struct packed {
      wt_cache_pkg::icache_in_t rtype;  // see definitions above
      logic [CVA6Cfg.ICACHE_LINE_WIDTH-1:0] data;  // full cache line width
      logic [CVA6Cfg.ICACHE_USER_LINE_WIDTH-1:0] user;  // user bits
      struct packed {
        logic                                      vld;  // invalidate only affected way
        logic                                      all;  // invalidate all ways
        logic [CVA6Cfg.ICACHE_INDEX_WIDTH-1:0]     idx;  // physical address to invalidate
        logic [CVA6Cfg.ICACHE_SET_ASSOC_WIDTH-1:0] way;  // way to invalidate
      } inv;  // invalidation vector
      logic [CVA6Cfg.MEM_TID_WIDTH-1:0] tid;  // threadi id (used as transaction id in Ariane)
    },

    // D$ data requests
    localparam type dcache_req_i_t = struct packed {
      logic [CVA6Cfg.DCACHE_INDEX_WIDTH-1:0] address_index;
      logic [CVA6Cfg.DCACHE_TAG_WIDTH-1:0]   address_tag;
      logic [CVA6Cfg.XLEN-1:0]               data_wdata;
      logic [CVA6Cfg.DCACHE_USER_WIDTH-1:0]  data_wuser;
      logic                                  data_req;
      logic                                  data_we;
      logic [(CVA6Cfg.XLEN/8)-1:0]           data_be;
      logic [1:0]                            data_size;
      logic [CVA6Cfg.DcacheIdWidth-1:0]      data_id;
      logic                                  kill_req;
      logic                                  tag_valid;
    },

    localparam type dcache_req_o_t = struct packed {
      logic                                 data_gnt;
      logic                                 data_rvalid;
      logic [CVA6Cfg.DcacheIdWidth-1:0]     data_rid;
      logic [CVA6Cfg.XLEN-1:0]              data_rdata;
      logic [CVA6Cfg.DCACHE_USER_WIDTH-1:0] data_ruser;
    },

    // AXI types
    parameter type axi_ar_chan_t = struct packed {
      logic [CVA6Cfg.AxiIdWidth-1:0]   id;
      logic [CVA6Cfg.AxiAddrWidth-1:0] addr;
      axi_pkg::len_t                   len;
      axi_pkg::size_t                  size;
      axi_pkg::burst_t                 burst;
      logic                            lock;
      axi_pkg::cache_t                 cache;
      axi_pkg::prot_t                  prot;
      axi_pkg::qos_t                   qos;
      axi_pkg::region_t                region;
      logic [CVA6Cfg.AxiUserWidth-1:0] user;
    },
    parameter type axi_aw_chan_t = struct packed {
      logic [CVA6Cfg.AxiIdWidth-1:0]   id;
      logic [CVA6Cfg.AxiAddrWidth-1:0] addr;
      axi_pkg::len_t                   len;
      axi_pkg::size_t                  size;
      axi_pkg::burst_t                 burst;
      logic                            lock;
      axi_pkg::cache_t                 cache;
      axi_pkg::prot_t                  prot;
      axi_pkg::qos_t                   qos;
      axi_pkg::region_t                region;
      axi_pkg::atop_t                  atop;
      logic [CVA6Cfg.AxiUserWidth-1:0] user;
    },
    parameter type axi_w_chan_t = struct packed {
      logic [CVA6Cfg.AxiDataWidth-1:0]     data;
      logic [(CVA6Cfg.AxiDataWidth/8)-1:0] strb;
      logic                                last;
      logic [CVA6Cfg.AxiUserWidth-1:0]     user;
    },
    parameter type b_chan_t = struct packed {
      logic [CVA6Cfg.AxiIdWidth-1:0]   id;
      axi_pkg::resp_t                  resp;
      logic [CVA6Cfg.AxiUserWidth-1:0] user;
    },
    parameter type r_chan_t = struct packed {
      logic [CVA6Cfg.AxiIdWidth-1:0]   id;
      logic [CVA6Cfg.AxiDataWidth-1:0] data;
      axi_pkg::resp_t                  resp;
      logic                            last;
      logic [CVA6Cfg.AxiUserWidth-1:0] user;
    },
    parameter type noc_req_t = struct packed {
      axi_aw_chan_t aw;
      logic         aw_valid;
      axi_w_chan_t  w;
      logic         w_valid;
      logic         b_ready;
      axi_ar_chan_t ar;
      logic         ar_valid;
      logic         r_ready;
    },
    parameter type noc_resp_t = struct packed {
      logic    aw_ready;
      logic    ar_ready;
      logic    w_ready;
      logic    b_valid;
      b_chan_t b;
      logic    r_valid;
      r_chan_t r;
    },
    //
    parameter type acc_cfg_t = logic,
    parameter acc_cfg_t AccCfg = '0
) (
    // Subsystem Clock - SUBSYSTEM
    input logic clk_i,
    // Asynchronous reset active low - SUBSYSTEM
    input logic rst_ni,
    // Reset boot address - SUBSYSTEM
    input logic [CVA6Cfg.VLEN-1:0] boot_addr_i,
    // Hard ID reflected as CSR - SUBSYSTEM
    input logic [CVA6Cfg.XLEN-1:0] hart_id_i,
    // Level sensitive (async) interrupts - SUBSYSTEM
    input logic [1:0] irq_i,
    // Inter-processor (async) interrupt - SUBSYSTEM
    input logic ipi_i,
    // Timer (async) interrupt - SUBSYSTEM
    input logic time_irq_i,
    // Debug (async) request - SUBSYSTEM
    input logic debug_req_i,
    // Probes to build RVFI, can be left open when not used - RVFI
    output rvfi_probes_t rvfi_probes_o,
	output wire         m_axi_ctrl_AWVALID,
	input  wire         m_axi_ctrl_AWREADY, //
	output wire [5:0]   m_axi_ctrl_AWID,
	output wire [63:0]  m_axi_ctrl_AWADDR,
	output wire [2:0]   m_axi_ctrl_AWSIZE,
	output wire [7:0]   m_axi_ctrl_AWLEN,
	output wire [1:0]   m_axi_ctrl_AWBURST,
	output wire         m_axi_ctrl_WVALID,
	input  wire         m_axi_ctrl_WREADY, //
	output wire [63:0]  m_axi_ctrl_WDATA,
	output wire [7:0]   m_axi_ctrl_WSTRB,
	output wire         m_axi_ctrl_WLAST,
	input  wire         m_axi_ctrl_BVALID, //
	output wire         m_axi_ctrl_BREADY,
	input  wire [5:0]   m_axi_ctrl_BID, //
	input  wire [1:0]   m_axi_ctrl_BRESP, //
	
	output wire         m_axi_ctrl_ARVALID,
	input  wire         m_axi_ctrl_ARREADY,//
	output wire [5:0]   m_axi_ctrl_ARID,
	output wire [63:0]  m_axi_ctrl_ARADDR,
	output wire [2:0]   m_axi_ctrl_ARSIZE,
	output wire [7:0]   m_axi_ctrl_ARLEN,
	output wire [1:0]   m_axi_ctrl_ARBURST,

    output wire [1:0]   m_axi_ctrl_ARPROT,
    output wire [1:0]   m_axi_ctrl_AWPROT,
	
	input  wire         m_axi_ctrl_RVALID, //
	output wire         m_axi_ctrl_RREADY,
	input  wire [5:0]   m_axi_ctrl_RID, //
	input  wire [63:0]  m_axi_ctrl_RDATA, //
	input  wire [1:0]   m_axi_ctrl_RRESP, //
	input  wire         m_axi_ctrl_RLAST, //

    output logic        EN_ctx_mem_access,
    output logic        ctx_mem_wr_en,
    output logic [31:0] ctx_mem_addr,
    output logic [31:0] ctx_mem_wr_data,

    input logic        ctx_mem_rd_resp_valid,
    input logic [31:0] ctx_mem_rd_data

);
noc_resp_t noc_resp;
noc_req_t noc_req;

assign noc_resp.aw_ready = m_axi_ctrl_AWREADY;
assign noc_resp.ar_ready = m_axi_ctrl_ARREADY;
assign noc_resp.w_ready = m_axi_ctrl_WREADY;
assign noc_resp.b_valid = m_axi_ctrl_BVALID;
assign noc_resp.b.id = m_axi_ctrl_BID;
assign noc_resp.b.resp = m_axi_ctrl_BRESP;
assign noc_resp.b.user = 0;
assign noc_resp.r_valid = m_axi_ctrl_RVALID;
assign noc_resp.r.id = m_axi_ctrl_RID;
assign noc_resp.r.data = m_axi_ctrl_RDATA;
assign noc_resp.r.resp = m_axi_ctrl_RRESP;
assign noc_resp.r.last = m_axi_ctrl_RLAST;

assign m_axi_ctrl_AWVALID =  noc_req.aw_valid;
assign m_axi_ctrl_AWID =  noc_req.aw.id;
assign m_axi_ctrl_AWADDR =  noc_req.aw.addr;
assign m_axi_ctrl_AWSIZE =  noc_req.aw.size;
assign m_axi_ctrl_AWLEN =  noc_req.aw.len;
assign m_axi_ctrl_AWBURST =  noc_req.aw.burst;
assign m_axi_ctrl_WVALID =  noc_req.w_valid;
assign m_axi_ctrl_WDATA =  noc_req.w.data;
assign m_axi_ctrl_WSTRB =  noc_req.w.strb;
assign m_axi_ctrl_WLAST =  noc_req.w.last;
assign m_axi_ctrl_BREADY =  noc_req.b_ready;
assign m_axi_ctrl_ARVALID =  noc_req.ar_valid;
assign m_axi_ctrl_ARID =  noc_req.ar.id;
assign m_axi_ctrl_ARADDR =  noc_req.ar.addr;
assign m_axi_ctrl_ARSIZE =  noc_req.ar.size;
assign m_axi_ctrl_ARLEN =  noc_req.ar.len;
assign m_axi_ctrl_ARBURST =  noc_req.ar.burst;
assign m_axi_ctrl_RREADY =  noc_req.r_ready;

assign m_axi_ctrl_ARPROT = 'b11;
assign m_axi_ctrl_AWPROT = 'b11;

// cva6 <-> ctx wiring
logic ctx_trap;
logic ctx_mret;

logic        ctx_inst_en;
logic  [2:0] ctx_inst_funct3;
logic [31:0] ctx_inst_rs1;
logic [31:0] ctx_inst_rs2;
logic [32:0] ctx_inst_rd;

//ctx
logic [31:0] ctx_mstatus;
logic [31:0] ctx_mepc;
logic [31:0] ctx_mcause;
logic        ctx_stall_mret;

logic         ctx_write_csrs;
logic  [31:0] ctx_mepc_rest;
logic  [31:0] ctx_mstatus_rest;

// rf access
logic        switch_bank;
logic [ 4:0] raddr_cold;
logic [31:0] rdata_cold;
logic [ 4:0] waddr_cold;
logic [31:0] wdata_cold;
logic        we_cold;

// write request separation
logic [36:0] reg_write_cold_u_to_c;
assign waddr_cold = reg_write_cold_u_to_c[36:32];
assign wdata_cold = reg_write_cold_u_to_c[31:0];

// memory access arbitration
logic RDY_ctx_mem_access;
logic [64:0] ctx_mem_access;

assign EN_ctx_mem_access = ~m_axi_ctrl_AWVALID & ~m_axi_ctrl_ARVALID & RDY_ctx_mem_access;
assign ctx_mem_addr      = ctx_mem_access[64:33];
assign ctx_mem_wr_data   = ctx_mem_access[32:1];
assign ctx_mem_wr_en     = ctx_mem_access[0];

// hot regs
logic [5:0] ctx_reg_hot_write_trace;

// Instantiate mkRTOSUnitSynth
mkRTOSUnitSynth u_mkRTOSUnitSynth (
    .CLK                        (clk_i),                      // Clock input
    .RST_N                      (rst_ni),                    // Reset input

    // Register Read Logic
    .reg_read_addr_cold         (raddr_cold), // reg_read_addr_cold
    .reg_read_data_cold_data    (rdata_cold), // reg_read_data_cold_data

    // Register Write Logic
    .EN_reg_write_cold          (we_cold), // EN_reg_write_cold
    .reg_write_cold             (reg_write_cold_u_to_c),    // reg_write_cold
    .RDY_reg_write_cold         (we_cold), // RDY_reg_write_cold

    // Cold Registers Logic
    .cold_regs_in               (928'b0),      // cold_regs_in

    // Hot Register Write Logic
    .reg_hot_write_trace_addrs   ({6'b0, ctx_reg_hot_write_trace}), // reg_hot_write_trace_addr

    // Memory Read Data Logic
    .mem_rd_data_d              (ctx_mem_rd_data),     // mem_rd_data_d
    .EN_mem_rd_data             (ctx_mem_rd_resp_valid),    // EN_mem_rd_data

    .mem_access                 (ctx_mem_access),
    .EN_mem_access              (EN_ctx_mem_access),
    .RDY_mem_access             (RDY_ctx_mem_access),

    // Mstatus and Mepc Logic
    .mstatus_out                (ctx_mstatus_rest),       // mstatus_out
    .mepc_out                   (ctx_mepc_rest),          // mepc_out

    // Bank Switching Logic
    .switch_bank_o              (switch_bank),     // switch_bank_o

    // Mret Logic
    .EN_mret                    (ctx_mret),           // EN_mret
    .mret                       (),              // mret
    .RDY_mret                   (ctx_stall_mret),          // RDY_mret

    // CSR Write Logic
    .write_csrs                 (ctx_write_csrs),        // write_csrs

    // Trap Logic
    .trap_mstatus               (ctx_mstatus),      // trap_mstatus
    .trap_mepc                  (ctx_mepc),         // trap_mepc
    .trap_mcause                (ctx_mcause),       // trap_mcause
    .EN_trap                    (ctx_trap),           // EN_trap
    .RDY_trap                   (),          // RDY_trap

    // Custom Instruction Logic
    .custom_inst_funct3         (ctx_inst_funct3),// custom_inst_funct3
    .custom_inst_id             (ctx_inst_rs1),    // custom_inst_id
    .custom_inst_prio           (ctx_inst_rs2),  // custom_inst_prio
    .EN_custom_inst             (ctx_inst_en),    // EN_custom_inst
    .custom_inst                (ctx_inst_rd),       // custom_inst
    .RDY_custom_inst            ()    // RDY_custom_inst
);

cva6 #(.CVA6Cfg ( CVA6Cfg )) cva6(
    .clk_i,
    .rst_ni,
    .boot_addr_i,
    .hart_id_i,
    .irq_i,
    .ipi_i,
    .time_irq_i,
    .debug_req_i,
    .cvxif_resp_i(113'b0),
    .cvxif_req_o(),
    .noc_resp_i(noc_resp),
    .noc_req_o(noc_req),
    .rvfi_probes_o(),

    .ctx_trap_o(ctx_trap),
    .ctx_mret_o(ctx_mret),

    .ctx_inst_funct3_o (ctx_inst_funct3),
    .ctx_inst_rs1_o    (ctx_inst_rs1),
    .ctx_inst_rs2_o    (ctx_inst_rs2),
    .ctx_inst_en_o     (ctx_inst_en),
    .ctx_inst_rd_i     (ctx_inst_rd[31:0]),

    //ctx
    .ctx_mstatus_o(ctx_mstatus),
    .ctx_mepc_o(ctx_mepc),
    .ctx_mcause_o(ctx_mcause),

    .switch_bank_i(switch_bank),
    .raddr_cold_i(raddr_cold),
    .rdata_cold_o(rdata_cold),
    .waddr_cold_i(waddr_cold),
    .wdata_cold_i(wdata_cold),
    .we_cold_i(we_cold),

    .ctx_stall_i(~ctx_stall_mret),

    .ctx_write_csrs_i(ctx_write_csrs),
    .ctx_mepc_i(ctx_mepc_rest),
    .ctx_mstatus_i(ctx_mstatus_rest),

    .ctx_reg_hot_write_trace_o(ctx_reg_hot_write_trace)
  );

endmodule
